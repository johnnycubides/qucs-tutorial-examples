* Qucs 0.0.24 /home/johnny/projects/qucs-tutorial-examples/examples/bjt/bjt1.sch
.INCLUDE "/tmp/.mount_qucs.ajpBTVx/usr/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"
* Qucs 0.0.24  /home/johnny/projects/qucs-tutorial-examples/examples/bjt/bjt1.sch
QT_2N2222_1 vout vb ve QMOD_T_2N2222_1 AREA=1.0 TEMP=26.85
.MODEL QMOD_T_2N2222_1 npn (Is=1e-14 Nf=1 Nr=1 Ikf=0.3 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=200 Br=3 Rbm=0 Irb=0 Rc=3 Re=1 Rb=10 Cje=2.5e-11 Vje=0.75 Mje=0.33 Cjc=8e-12 Vjc=0.75 Mjc=0.33 Xcjc=1 Cjs=0 Vjs=0.75 Mjs=0 Fc=0.5 Tf=4e-10 Xtf=3 Vtf=0 Itf=2 Tr=1e-07 Kf=0 Af=1 Ptf=0 Xtb=0 Xti=3 Eg=1.11 Tnom=26.85 )
V1 vcc 0 DC 15
R1 vb vcc  10K
R2 0 vb  2K
R4 vout vcc  1K
R3 0 ve  100
EPr1 Pr1 0 vout 0 1.0
RPr1Pr1 Pr1 0 1E8
RPr1vout vout 0 1E8
EPr2 Pr2 0 ve 0 1.0
RPr2Pr2 Pr2 0 1E8
RPr2ve ve 0 1E8
.control
echo "" > spice4qucs.cir.noise
echo "" > spice4qucs.cir.pz
tran 9.09091e-05 0.001 0 
write bjt1_tran.txt v(Pr1) v(Pr2) v(vb) v(vcc) v(ve) v(vout) 
destroy all
reset

exit
.endc
.END
